spi_PLL_inst : spi_PLL PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
